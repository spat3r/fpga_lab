module hdmi_fir_IP #(
    //TODO: add some parameters
) (
    //TODO: add some ports
);
    // TODO: Instanciate fir_axi_if.sv


    // TODO: Instanuciate hdmi_top.sv


    // TODO: reading histogram bins


    // TODO: writing fir parameters

    // TODO: szerintem az axi regiszterek itt legyenek implementálva és az almodulok csak hozzáférnek vezetékeken keresztül
                // biztosan egy vezetékezési kín lesz de nem tudom hogy lehet optimálisan megoldani
endmodule