module fir_axi_if #(
    //TODO: add parameters
) (
    //TODO: add ports
);
// TODO: Kell készíteni egy AXI interfész modult (nem tudom fel lehet e használni a fluid leveleset.)
    //TODO: implement fsm

    //TODO implement fir writing, bin reading
endmodule