module fir_axi_if #(
    //TODO: add parameters
) (
    //TODO: add ports
);
    //TODO: implement fsm

    //TODO implement fir writing, bin reading
endmodule